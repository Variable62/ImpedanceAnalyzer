module PhaseCounter (
    input       wire        Clk48,
    input       wire        ExtResetn,

);
    
endmodule